// Copyright 2023 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Yvan Tortorella <yvan.tortorella@unibo.it>
//

timeunit 1ps; timeprecision 1ps;

import hci_package::*;

module redmule_tb

  import redmule_pkg::*;
#(
  parameter TCP = 1.0ns, // clock period, 1 GHz clock
  parameter TA  = 0.2ns, // application time
  parameter TT  = 0.8ns,  // test time
  parameter logic UseXif = 1'b0,
  parameter real  PROB_STALL = 0,
  parameter logic mx_enable = 1'b1
)(
  input logic clk_i,
  input logic rst_ni,
  input logic fetch_enable_i
);

  // parameters
  // MX test vector storage for data - NO LONGER NEEDED: data compiled from C headers
  // logic [15:0] mx_x_data_mem [0:511];  // 512 16-bit words (1024 FP8 values packed)
  // logic [15:0] mx_w_data_mem [0:511];  // 512 16-bit words (1024 FP8 values packed)

  localparam int unsigned NC = 1;
  localparam int unsigned ID = 10;
  localparam int unsigned DW = redmule_pkg::DATA_W;
  localparam int unsigned MP = DW/32;
  localparam int unsigned MEMORY_SIZE = 192*1024;
  localparam int unsigned STACK_MEMORY_SIZE = 192*1024;
  localparam int unsigned PULP_XPULP = 1;
  localparam int unsigned FPU = 0;
  localparam int unsigned PULP_ZFINX = 0;
  localparam logic [31:0] BASE_ADDR = 32'h1c000000;
  localparam logic [31:0] DUMMY_DMEM_BASE = 32'h1c010000;
  localparam logic [31:0] X_EXP_BASE_ADDR = BASE_ADDR + 32'h0002_0000;
  localparam logic [31:0] W_EXP_BASE_ADDR = BASE_ADDR + 32'h0002_1000;
  localparam int unsigned X_EXP_MEM_OFFSET = (X_EXP_BASE_ADDR - DUMMY_DMEM_BASE) >> 2;
  localparam int unsigned W_EXP_MEM_OFFSET = (W_EXP_BASE_ADDR - DUMMY_DMEM_BASE) >> 2;
  localparam logic [31:0] HWPE_ADDR_BASE_BIT = 20;
  localparam bit          USE_ECC = 0;
  localparam int unsigned EW = (USE_ECC) ? 72 : DEFAULT_EW;
  localparam redmule_pkg::core_type_e CoreType = UseXif ? redmule_pkg::CV32X
                                                        : redmule_pkg::CV32P;

  localparam hci_package::hci_size_parameter_t HciRedmuleSize = '{
    DW:  DW,
    AW:  hci_package::DEFAULT_AW,
    BW:  hci_package::DEFAULT_BW,
    UW:  hci_package::DEFAULT_UW,
    IW:  hci_package::DEFAULT_IW,
    EW:  EW,
    EHW: hci_package::DEFAULT_EHW,
    default: '0
  };


  // global signals
  string stim_instr, stim_data, stack_init;
  string x_exp_file, w_exp_file;
  string mx_dir_resolved; // Directory for MX vectors, derived from stim_data
  logic test_mode;
  logic [31:0] core_boot_addr;
  logic redmule_busy;
  logic core_sleep;
  int errors;
  integer f_engine_x, f_engine_w, f_engine_z;
  integer f_dec_fp16, f_dec_exp, f_dec_target;

  task automatic load_exponent_file(string path, int base_word_offset);
    int fd;
    int idx;
    int word_val;
    fd = $fopen(path, "r");
    if (!fd) begin
      $fatal(1, "[TB] Failed to open exponent file %s", path);
    end
    idx = 0;
    // Compact format: read 32-bit words directly (no padding)
    // Each line in the file is one 32-bit word in hex
    while (!$feof(fd)) begin
      if ($fscanf(fd, "%h\n", word_val) != 1) begin
        break;
      end
      // Store directly as 32-bit word - streamer will read 512-bit beats (16 words)
      i_dummy_dmemory.memory[base_word_offset + idx] = word_val;
      idx++;
    end
    $fclose(fd);
    $display("[TB] Loaded %0d exponent words from %s", idx, path);
  endtask

  // ---------------------------------------------------------------------------
  // Performance counters
  // ---------------------------------------------------------------------------
  bit perf_enable;
  logic perf_active;
  logic perf_seen_busy; // Track if we've seen busy_o high during this measurement
  longint unsigned perf_total_cycles;
  longint unsigned perf_busy_cycles;
  longint unsigned perf_encoder_blocks;
  longint unsigned perf_decoder_blocks;

  // Optional MX debug dumping (enabled with +MX_DEBUG_DUMP)
  bit mx_debug_dump;
  integer mx_debug_fd;
  initial begin
    mx_debug_dump = 1'b1;
    mx_debug_fd   = $fopen("mx_debug.log", "w");
    if (mx_debug_fd == 0) begin
      $display("[TB][MXDBG] Failed to open mx_debug.log, disabling dump");
      mx_debug_dump = 1'b0;
    end else begin
      $display("[TB][MXDBG] Logging MX slot/decoder activity to mx_debug.log");
      $fdisplay(mx_debug_fd,
                "time,stage,target,data,exp");
    end
  end

  final begin
    if (mx_debug_dump) begin
      $fclose(mx_debug_fd);
    end
    if (f_engine_x) $fclose(f_engine_x);
    if (f_engine_w) $fclose(f_engine_w);
    if (f_engine_z) $fclose(f_engine_z);
    if (f_dec_fp16) $fclose(f_dec_fp16);
    if (f_dec_exp) $fclose(f_dec_exp);
    if (f_dec_target) $fclose(f_dec_target);
    $writememh("y_oup_dump.mem", redmule_tb.i_dummy_dmemory.memory);
  end

  initial begin
    if (!$value$plusargs("PERF_ENABLE=%0d", perf_enable)) begin
      perf_enable = 1'b1;
    end
  end

  // Engine/decoder dump files
  initial begin
    f_engine_x = $fopen("engine_x_inputs.txt", "w");
    if (f_engine_x == 0) begin
      $fatal(1, "[TB] Failed to open engine_x_inputs.txt");
    end
    f_engine_w = $fopen("engine_w_inputs.txt", "w");
    if (f_engine_w == 0) begin
      $fatal(1, "[TB] Failed to open engine_w_inputs.txt");
    end
    f_engine_z = $fopen("engine_z_outputs.txt", "w");
    if (f_engine_z == 0) begin
      $fatal(1, "[TB] Failed to open engine_z_outputs.txt");
    end
    f_dec_fp16 = $fopen("mx_decoder_fp16_outputs.txt", "w");
    if (f_dec_fp16 == 0) begin
      $fatal(1, "[TB] Failed to open mx_decoder_fp16_outputs.txt");
    end
    f_dec_exp = $fopen("mx_decoder_exponents.txt", "w");
    if (f_dec_exp == 0) begin
      $fatal(1, "[TB] Failed to open mx_decoder_exponents.txt");
    end
    f_dec_target = $fopen("mx_decoder_targets.txt", "w");
    if (f_dec_target == 0) begin
      $fatal(1, "[TB] Failed to open mx_decoder_targets.txt");
    end
  end

  // Performance counters measure full accelerator execution including MX encoding/decoding
  // Start: busy_o rises OR first TCDM request OR first MX encoder/decoder activity
  // Stop: Timeout after last activity (busy, TCDM, or MX encoder/decoder)

  logic accel_active; // Combined activity signal
  int idle_count;     // Count idle cycles for timeout
  localparam int IDLE_TIMEOUT = 10; // Cycles of inactivity before stopping measurement

  // Debug counters for stream completions
  int x_stream_done_count;
  int w_stream_done_count;
  int z_stream_done_count;

  assign accel_active = i_dut.i_redmule_top.busy_o ||
                        redmule_tcdm.req ||
                        (i_dut.i_redmule_top.mx_val_valid && i_dut.i_redmule_top.mx_val_ready) ||
                        (i_dut.i_redmule_top.mx_dec_fp16_valid && i_dut.i_redmule_top.mx_dec_fp16_ready);

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      perf_active         <= 1'b0;
      perf_seen_busy      <= 1'b0;
      perf_total_cycles   <= '0;
      perf_busy_cycles    <= '0;
      perf_encoder_blocks <= '0;
      perf_decoder_blocks <= '0;
      idle_count          <= 0;
      x_stream_done_count <= 0;
      w_stream_done_count <= 0;
      z_stream_done_count <= 0;
    end else begin
      if (perf_enable) begin
        // Track stream completions using hci_streamer_flags_t.done field
        if (i_dut.i_redmule_top.flgs_streamer.x_stream_source_flags.done)
          x_stream_done_count <= x_stream_done_count + 1;
        if (i_dut.i_redmule_top.flgs_streamer.w_stream_source_flags.done)
          w_stream_done_count <= w_stream_done_count + 1;
        if (i_dut.i_redmule_top.flgs_streamer.z_stream_sink_flags.done)
          z_stream_done_count <= z_stream_done_count + 1;

        if (!perf_active) begin
          // Start measurement on first activity after fetch_enable
          if (fetch_enable_i && accel_active) begin
            perf_active <= 1'b1;
            idle_count <= 0;
          end
        end else begin
          // Measurement active: track cycles and activity
          perf_total_cycles <= perf_total_cycles + 1;

          if (i_dut.i_redmule_top.busy_o) begin
            perf_busy_cycles <= perf_busy_cycles + 1;
            perf_seen_busy <= 1'b1;
          end

          if (i_dut.i_redmule_top.mx_val_valid && i_dut.i_redmule_top.mx_val_ready) begin
            perf_encoder_blocks <= perf_encoder_blocks + 1;
          end

          if (i_dut.i_redmule_top.mx_dec_fp16_valid && i_dut.i_redmule_top.mx_dec_fp16_ready) begin
            perf_decoder_blocks <= perf_decoder_blocks + 1;
            if (f_dec_fp16) begin
              // mx_dec_fp16_data is a flat vector (NUM_LANES*BITW), so slice per lane
              for (int lane = 0; lane < ARRAY_WIDTH; lane++) begin
                $fwrite(f_dec_fp16,
                        "%04h ",
                        i_dut.i_redmule_top.mx_dec_fp16_data[lane*BITW +: BITW]);
              end
              $fwrite(f_dec_fp16, "\n");
            end
            if (f_dec_target) begin
              if (i_dut.i_redmule_top.target_is_x) begin
                $fwrite(f_dec_target, "X\n");
              end else if (i_dut.i_redmule_top.target_is_w) begin
                $fwrite(f_dec_target, "W\n");
              end else begin
                $fwrite(f_dec_target, "-\n");
              end
            end
          end

          // Timeout logic: stop after IDLE_TIMEOUT cycles of no activity
          if (accel_active) begin
            idle_count <= 0;
          end else begin
            idle_count <= idle_count + 1;
            if (idle_count >= IDLE_TIMEOUT && perf_seen_busy) begin
              perf_active <= 1'b0;
              perf_seen_busy <= 1'b0;
              idle_count <= 0;
            end
          end
        end
      end

      if (perf_active && core_sleep && (errors != -1)) begin
        perf_active <= 1'b0;
      end
    end
  end
  logic scan_cg_en;

  // Log MX decoder exponents whenever the decoder accepts a new block
  always @(posedge clk_i) begin
    if (f_dec_exp &&
        i_dut.i_redmule_top.mx_dec_exp_valid &&
        i_dut.i_redmule_top.mx_dec_exp_ready) begin
      $fwrite(f_dec_exp, "%0h\n", i_dut.i_redmule_top.mx_dec_exp_data);
    end
  end

  // Helper: get directory name from path
  function automatic string dirname(input string path);
    int i;
    dirname = path;
    // find last '/'
    for (i = path.len()-1; i >= 0; i--) begin
      if (path.getc(i) == "/") begin
        dirname = path.substr(0, i-1);
        return dirname;
      end
    end
    // no slash -> current dir
    dirname = ".";
  endfunction

  hwpe_stream_intf_tcdm instr[0:0]  (.clk(clk_i));
  hwpe_stream_intf_tcdm stack[0:0]  (.clk(clk_i));
  hwpe_stream_intf_tcdm tcdm [MP:0] (.clk(clk_i));
  
  // MX exponent stream interface (encoder output)
  hwpe_stream_intf_stream #(.DATA_WIDTH(32)) mx_exp_stream (.clk(clk_i));

  // Drive ready to always accept encoder exponent outputs
  assign mx_exp_stream.ready = 1'b1;
  
    logic [NC-1:0][1:0]  evt;
  logic [MP-1:0]       tcdm_gnt;
  logic [MP-1:0][31:0] tcdm_r_data;
  logic [MP-1:0]       tcdm_r_valid;

  typedef struct packed {
    logic        req;
    logic [31:0] addr;
  } core_inst_req_t;

  typedef struct packed {
    logic        gnt;
    logic        valid;
    logic [31:0] data;
  } core_inst_rsp_t;

  typedef struct packed {
    logic req;
    logic we;
    logic [3:0] be;
    logic [31:0] addr;
    logic [31:0] data;
  } core_data_req_t;

  typedef struct packed {
    logic gnt;
    logic valid;
    logic [31:0] data;
  } core_data_rsp_t;

  hci_core_intf #(.DW(DW)) redmule_tcdm (.clk(clk_i));

  core_inst_req_t core_inst_req;
  core_inst_rsp_t core_inst_rsp;

  core_data_req_t core_data_req;
  core_data_rsp_t core_data_rsp;

  always_comb begin : bind_instrs
    instr[0].req  = core_inst_req.req;
    instr[0].add  = core_inst_req.addr;
    instr[0].wen  = 1'b1;
    instr[0].be   = '0;
    instr[0].data = '0;
    core_inst_rsp.gnt   = instr[0].gnt;
    core_inst_rsp.valid = instr[0].r_valid;
    core_inst_rsp.data  = instr[0].r_data;
  end

  always_comb begin : bind_stack
    stack[0].req  = core_data_req.req & (core_data_req.addr[31:16] == 16'h1c04) &
                    ~core_data_req.addr[HWPE_ADDR_BASE_BIT];
    stack[0].add  = core_data_req.addr;
    stack[0].wen  = ~core_data_req.we;
    stack[0].be   = core_data_req.be;
    stack[0].data = core_data_req.data;
  end

  logic other_r_valid;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (~rst_ni)
      other_r_valid <= '0;
    else
      other_r_valid <= core_data_req.req & (core_data_req.addr[31:24] == 8'h80);
  end

  for(genvar ii=0; ii<MP; ii++) begin : tcdm_binding
    assign tcdm[ii].req  = redmule_tcdm.req;
    assign tcdm[ii].add  = redmule_tcdm.add + ii*4;
    assign tcdm[ii].wen  = redmule_tcdm.wen;
    assign tcdm[ii].be   = redmule_tcdm.be[(ii+1)*4-1:ii*4];
    assign tcdm_gnt[ii]     = tcdm[ii].gnt;
    assign tcdm_r_valid[ii] = tcdm[ii].r_valid;
    assign tcdm_r_data[ii]  = tcdm[ii].r_data;
  end
  assign redmule_tcdm.gnt     = &tcdm_gnt;
  assign redmule_tcdm.r_data  = { >> {tcdm_r_data} };
  assign redmule_tcdm.r_valid = &tcdm_r_valid;
  assign redmule_tcdm.r_id    = '0;
  assign redmule_tcdm.r_opc   = '0;
  assign redmule_tcdm.r_user  = '0;

  if (USE_ECC) begin : gen_ecc
    logic [EW-1:0] tcdm_r_ecc;
    // RESPONSE PHASE ENCODING
    logic [MP-1:0][38:0] tcdm_r_data_enc;
    for(genvar ii=0; ii<MP; ii++) begin : gen_rdata_encoders
      hsiao_ecc_enc #(
        .DataWidth ( 32 )
      ) i_r_data_enc (
        .in  (tcdm_r_data[ii]),
        .out (tcdm_r_data_enc[ii])
      );
      assign tcdm_r_ecc[(ii+1)*7-1:ii*7] = tcdm_r_data_enc[ii][38:32];
    end
    assign tcdm_r_ecc[EW-1:(7*MP)] = '0;
    assign redmule_tcdm.r_ecc  = tcdm_r_ecc;

    // REQUEST PHASE DECODING
    for(genvar ii=0; ii<MP; ii++) begin : gen_data_decoders
      hsiao_ecc_dec #(
        .DataWidth ( 32 )
      ) i_data_dec (
        .in         ( { redmule_tcdm.ecc[(ii+1)*7-1+9:ii*7+9], redmule_tcdm.data[(ii+1)*32-1:ii*32] } ),
        .out        ( tcdm[ii].data ),
        .syndrome_o ( ),
        .err_o      ( )
      );
    end

    // FixMe: How should we drive these?
    // assign redmule_tcdm.egnt = '1;
    // assign redmule_tcdm.r_evalid = '0;

  end else begin: gen_no_ecc
    for(genvar ii=0; ii<MP; ii++)
      assign tcdm[ii].data = redmule_tcdm.data[(ii+1)*32-1:ii*32];

    assign redmule_tcdm.r_ecc = '0;
    assign redmule_tcdm.egnt = '1;
    assign redmule_tcdm.r_evalid = '0;
  end

  assign tcdm[MP].req  = core_data_req.req &
                         (core_data_req.addr[31:24] != '0) &
                         (core_data_req.addr[31:24] != 8'h80) &
                         ~core_data_req.addr[HWPE_ADDR_BASE_BIT];
  assign tcdm[MP].add  = core_data_req.addr;
  assign tcdm[MP].wen  = ~core_data_req.we;
  assign tcdm[MP].be   = core_data_req.be;
  assign tcdm[MP].data = core_data_req.data;

  assign core_data_rsp.gnt = stack[0].req ?
                             stack[0].gnt : tcdm[MP].req ?
                                            tcdm[MP].gnt : '1;

  assign core_data_rsp.data = stack[0].r_valid ? stack[0].r_data  :
                                                 tcdm[MP].r_valid ? tcdm[MP].r_data : '0;
  assign core_data_rsp.valid = stack[0].r_valid |
                               tcdm[MP].r_valid |
                               other_r_valid    ;

  tb_dummy_memory  #(
    .MP             ( MP + 1        ),
    .MEMORY_SIZE    ( MEMORY_SIZE   ),
    .BASE_ADDR      ( 32'h1c010000  ),
    .PROB_STALL     ( PROB_STALL    ),
    .TCP            ( TCP           ),
    .TA             ( TA            ),
    .TT             ( TT            )
  ) i_dummy_dmemory (
    .clk_i          ( clk_i         ),
    .rst_ni         ( rst_ni        ),
    .clk_delayed_i  ( '0            ),
    .randomize_i    ( 1'b0          ),
    .enable_i       ( 1'b1          ),
    .stallable_i    ( 1'b1          ),
    .tcdm           ( tcdm          )
  );

  tb_dummy_memory  #(
    .MP             ( 1           ),
    .MEMORY_SIZE    ( MEMORY_SIZE ),
    .BASE_ADDR      ( BASE_ADDR   ),
    .PROB_STALL     ( 0           ),
    .TCP            ( TCP         ),
    .TA             ( TA          ),
    .TT             ( TT          )
  ) i_dummy_imemory (
    .clk_i          ( clk_i       ),
    .rst_ni         ( rst_ni      ),
    .clk_delayed_i  ( '0          ),
    .randomize_i    ( 1'b0        ),
    .enable_i       ( 1'b1        ),
    .stallable_i    ( 1'b0        ),
    .tcdm           ( instr       )
  );

  tb_dummy_memory       #(
    .MP                  ( 1                 ),
    .MEMORY_SIZE         ( STACK_MEMORY_SIZE ),
    .BASE_ADDR           ( BASE_ADDR         ),
    .PROB_STALL          ( 0                 ),
    .TCP                 ( TCP               ),
    .TA                  ( TA                ),
    .TT                  ( TT                )
  ) i_dummy_stack_memory (
    .clk_i               ( clk_i             ),
    .rst_ni              ( rst_ni            ),
    .clk_delayed_i       ( '0                ),
    .randomize_i         ( 1'b0              ),
    .enable_i            ( 1'b1              ),
    .stallable_i         ( 1'b0              ),
    .tcdm                ( stack             )
  );

`ifdef TARGET_VERILATOR
  assign scan_cg_en = UseXif ? 1'b1 : 1'b0;
`else
  assign scan_cg_en = 1'b0;
`endif
  redmule_complex #(
    .CoreType           ( CoreType            ), // CV32E40P, CV32E40X, IBEX, SNITCH, CVA6
    .ID_WIDTH           ( ID                  ),
    .N_CORES            ( NC                  ),
    .NumIrqs            ( 1                   ),
    .AddrWidth          ( 32                  ),
    .HciRedmuleSize     ( HciRedmuleSize      ),
    .core_data_req_t    ( core_data_req_t     ),
    .core_data_rsp_t    ( core_data_rsp_t     ),
    .core_inst_req_t    ( core_inst_req_t     ),
    .core_inst_rsp_t    ( core_inst_rsp_t     )
  ) i_dut               (
    .clk_i              ( clk_i            ),
    .rst_ni             ( rst_ni           ),
    .test_mode_i        ( test_mode        ),
    .fetch_enable_i     ( fetch_enable_i   ),
    .scan_cg_en_i       ( scan_cg_en       ),
    .redmule_clk_en_i   ( 1'b1             ),
    .boot_addr_i        ( core_boot_addr   ),
    .irq_i              ( '0               ),
    .irq_id_o           (                  ),
    .irq_ack_o          (                  ),
    .core_sleep_o       ( core_sleep       ),
    .core_inst_rsp_i    ( core_inst_rsp    ),
    .core_inst_req_o    ( core_inst_req    ),
    .core_data_rsp_i    ( core_data_rsp    ),
    .core_data_req_o    ( core_data_req    ),
    .tcdm               ( redmule_tcdm     ),
    .mx_exp_stream      ( mx_exp_stream    )
  );

  integer f_x, f_W, f_y, f_tau;
  integer f_engine_x, f_engine_w, f_engine_z;
  integer f_dec_fp16, f_dec_exp, f_dec_target;
  logic start;
  logic x_buf_read_q, w_buf_read_q;


  always_ff @(posedge clk_i)
  begin
    if((core_data_req.addr == 32'h80000000) &&
       (core_data_req.we & core_data_req.req == 1'b1)) begin
      errors = core_data_req.data;
    end
    if((core_data_req.addr == 32'h80000004 ) &&
       (core_data_req.we & core_data_req.req == 1'b1)) begin
      $write("%c", core_data_req.data);
    end
  end

  // Track buffer read strobes (one-cycle delayed output valid)
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      x_buf_read_q <= 1'b0;
      w_buf_read_q <= 1'b0;
    end else begin
      x_buf_read_q <= i_dut.i_redmule_top.x_buffer_ctrl.h_shift;
      w_buf_read_q <= i_dut.i_redmule_top.w_buffer_ctrl.shift;
    end
  end

  // MX debug dump: capture slot buffer and decoder activity when enabled
  always_ff @(posedge clk_i) begin
    if (mx_debug_dump) begin
      automatic string target_str;
      logic slot_fire_x, slot_fire_w;
      logic x_mux_push, w_mux_push;
      logic x_fifo_pop, w_fifo_pop;
      slot_fire_x = i_dut.i_redmule_top.consume_x_slot &&
                    i_dut.i_redmule_top.i_mx_slot_buffer.x_slot_valid_o &&
                    i_dut.i_redmule_top.i_mx_slot_buffer.x_slot_exp_valid_o;
      slot_fire_w = i_dut.i_redmule_top.consume_w_slot &&
                    i_dut.i_redmule_top.i_mx_slot_buffer.w_slot_valid_o &&
                    i_dut.i_redmule_top.i_mx_slot_buffer.w_slot_exp_valid_o;
      x_mux_push = i_dut.i_redmule_top.x_buffer_muxed.valid &&
                   i_dut.i_redmule_top.x_buffer_muxed.ready;
      w_mux_push = i_dut.i_redmule_top.w_buffer_muxed.valid &&
                   i_dut.i_redmule_top.w_buffer_muxed.ready;
      x_fifo_pop = i_dut.i_redmule_top.x_buffer_fifo.valid &&
                   i_dut.i_redmule_top.x_buffer_fifo.ready;
      w_fifo_pop = i_dut.i_redmule_top.w_buffer_fifo.valid &&
                   i_dut.i_redmule_top.w_buffer_fifo.ready;

      if (slot_fire_x) begin
        $display("[TB][MXDBG][%0t] SLOT_X data=%h exp=%h",
                 $time,
                 i_dut.i_redmule_top.i_mx_slot_buffer.x_slot_data_o,
                 i_dut.i_redmule_top.i_mx_slot_buffer.x_slot_exp_o);
        if (mx_debug_fd)
          $fdisplay(mx_debug_fd,
                    "%0t,SLOT,X,%h,%h",
                    $time,
                    i_dut.i_redmule_top.i_mx_slot_buffer.x_slot_data_o,
                    i_dut.i_redmule_top.i_mx_slot_buffer.x_slot_exp_o);
      end

      if (slot_fire_w) begin
        $display("[TB][MXDBG][%0t] SLOT_W data=%h exp=%h",
                 $time,
                 i_dut.i_redmule_top.i_mx_slot_buffer.w_slot_data_o,
                 i_dut.i_redmule_top.i_mx_slot_buffer.w_slot_exp_o);
        if (mx_debug_fd)
          $fdisplay(mx_debug_fd,
                    "%0t,SLOT,W,%h,%h",
                    $time,
                    i_dut.i_redmule_top.i_mx_slot_buffer.w_slot_data_o,
                    i_dut.i_redmule_top.i_mx_slot_buffer.w_slot_exp_o);
      end

      if (x_mux_push) begin
        $display("[TB][MXDBG][%0t] XBUF data=%h",
                 $time,
                 i_dut.i_redmule_top.x_buffer_muxed.data);
        if (mx_debug_fd)
          $fdisplay(mx_debug_fd,
                    "%0t,XBUF,%s,%h,%s",
                    $time,
                    i_dut.i_redmule_top.target_is_x ? "X" : "?",
                    i_dut.i_redmule_top.x_buffer_muxed.data,
                    "-");
      end

      if (w_mux_push) begin
        $display("[TB][MXDBG][%0t] WBUF data=%h",
                 $time,
                 i_dut.i_redmule_top.w_buffer_muxed.data);
        if (mx_debug_fd)
          $fdisplay(mx_debug_fd,
                    "%0t,WBUF,%s,%h,%s",
                    $time,
                    i_dut.i_redmule_top.target_is_w ? "W" : "?",
                    i_dut.i_redmule_top.w_buffer_muxed.data,
                    "-");
      end

      if (x_fifo_pop) begin
        $display("[TB][MXDBG][%0t] XFIFO data=%h",
                 $time,
                 i_dut.i_redmule_top.x_buffer_fifo.data);
        if (mx_debug_fd)
          $fdisplay(mx_debug_fd,
                    "%0t,XFIFO,X,%h,%s",
                    $time,
                    i_dut.i_redmule_top.x_buffer_fifo.data,
                    "-");
      end

      if (w_fifo_pop) begin
        $display("[TB][MXDBG][%0t] WFIFO data=%h",
                 $time,
                 i_dut.i_redmule_top.w_buffer_fifo.data);
        if (mx_debug_fd)
          $fdisplay(mx_debug_fd,
                    "%0t,WFIFO,W,%h,%s",
                    $time,
                    i_dut.i_redmule_top.w_buffer_fifo.data,
                    "-");
      end

      if (x_buf_read_q) begin
        $display("[TB][MXDBG][%0t] XBUFQ row=%0d data=%h",
                 $time,
                 i_dut.i_redmule_top.i_x_buffer.h_index_r,
                 i_dut.i_redmule_top.x_buffer_q);
        if (mx_debug_fd)
          $fdisplay(mx_debug_fd,
                    "%0t,XBUFQ,X,%h,%s",
                    $time,
                    i_dut.i_redmule_top.x_buffer_q,
                    "-");
        if (f_engine_x) begin
          for (int w_idx = 0; w_idx < ARRAY_WIDTH; w_idx++) begin
            for (int h_idx = 0; h_idx < ARRAY_HEIGHT; h_idx++) begin
              $fwrite(f_engine_x, "%04h ",
                      i_dut.i_redmule_top.x_buffer_q[w_idx][h_idx]);
            end
          end
          $fwrite(f_engine_x, "\n");
        end
      end

      if (w_buf_read_q) begin
        $display("[TB][MXDBG][%0t] WBUFQ data=%h",
                 $time,
                 i_dut.i_redmule_top.w_buffer_q);
        if (mx_debug_fd)
          $fdisplay(mx_debug_fd,
                    "%0t,WBUFQ,W,%h,%s",
                    $time,
                    i_dut.i_redmule_top.w_buffer_q,
                    "-");
        if (f_engine_w) begin
          for (int h_idx = 0; h_idx < ARRAY_HEIGHT; h_idx++) begin
            $fwrite(f_engine_w, "%04h ",
                    i_dut.i_redmule_top.w_buffer_q[h_idx]);
          end
          $fwrite(f_engine_w, "\n");
        end
      end

      if (i_dut.i_redmule_top.fifo_valid &&
          i_dut.i_redmule_top.fifo_pop) begin
        if (f_engine_z) begin
          for (int lane = 0; lane < ARRAY_WIDTH; lane++) begin
            $fwrite(f_engine_z, "%04h ",
                    i_dut.i_redmule_top.fifo_data_out[lane*BITW +: BITW]);
          end
          $fwrite(f_engine_z, "\n");
        end
      end

      if (i_dut.i_redmule_top.mx_dec_fp16_valid &&
          i_dut.i_redmule_top.mx_dec_fp16_ready) begin
        target_str = i_dut.i_redmule_top.target_is_x ? "X" :
                     i_dut.i_redmule_top.target_is_w ? "W" : "NONE";
        $display("[TB][MXDBG][%0t] DEC_%s data=%h",
                 $time,
                 target_str,
                 i_dut.i_redmule_top.mx_dec_fp16_data);
        if (mx_debug_fd)
          $fdisplay(mx_debug_fd,
                    "%0t,DEC,%s,%h,%s",
                    $time,
                    target_str,
                    i_dut.i_redmule_top.mx_dec_fp16_data,
                    "-");
      end
    end
  end

  initial begin
    integer id;
    int cnt_rd, cnt_wr;

    errors = -1;
    if (!$value$plusargs("STIM_INSTR=%s", stim_instr)) stim_instr = "";
    if (!$value$plusargs("STIM_DATA=%s", stim_data)) stim_data = "";
    if (!$value$plusargs("STACK_INIT=%s", stack_init)) stack_init = "";
    if (!$value$plusargs("X_EXP_FILE=%s", x_exp_file)) x_exp_file = "";
    if (!$value$plusargs("W_EXP_FILE=%s", w_exp_file)) w_exp_file = "";
    $display("Please find STIM_INSTR loaded from %s", stim_instr);
    $display("Please find STIM_DATA loaded from %s", stim_data);
    $display("Please find STACK_INIT loaded from %s", stack_init);

    // MX: derive exponent file paths from stim_data
    if (mx_enable) begin
      mx_dir_resolved = dirname(stim_data);
      $display("[TB] MX dir derived from STIM_DATA: %s", mx_dir_resolved);
      $display("[TB] FW is responsible for loading MX exponent tables");
    end

    test_mode = 1'b0;
    core_boot_addr = 32'h1C000084;

    // Load instruction and data memory
    $readmemh(stim_instr, redmule_tb.i_dummy_imemory.memory);
    $readmemh(stim_data,  redmule_tb.i_dummy_dmemory.memory);
    $readmemh(stack_init, redmule_tb.i_dummy_stack_memory.memory);
    // Firmware now loads MX exponent tables; no preload here
    // End: WFI + returned != -1 signals end-of-computation
    while(~core_sleep || errors==-1) begin
      // Feed MX data to X and W buffers if enabled
      if (mx_enable) begin
        // Example: drive X and W buffer inputs from test vectors
        // (Replace with actual buffer interface as needed)
        // x_buffer_data_in = mx_x_data_mem[mx_x_data_idx];
        // w_buffer_data_in = mx_w_data_mem[mx_w_data_idx];
      end
      @(posedge clk_i);
    end
    cnt_rd = redmule_tb.i_dummy_dmemory.cnt_rd[0] +
             redmule_tb.i_dummy_dmemory.cnt_rd[1] +
             redmule_tb.i_dummy_dmemory.cnt_rd[2] +
             redmule_tb.i_dummy_dmemory.cnt_rd[3] +
             redmule_tb.i_dummy_dmemory.cnt_rd[4] +
             redmule_tb.i_dummy_dmemory.cnt_rd[5] +
             redmule_tb.i_dummy_dmemory.cnt_rd[6] +
             redmule_tb.i_dummy_dmemory.cnt_rd[7] +
             redmule_tb.i_dummy_dmemory.cnt_rd[8];

    cnt_wr = redmule_tb.i_dummy_dmemory.cnt_wr[0] +
             redmule_tb.i_dummy_dmemory.cnt_wr[1] +
             redmule_tb.i_dummy_dmemory.cnt_wr[2] +
             redmule_tb.i_dummy_dmemory.cnt_wr[3] +
             redmule_tb.i_dummy_dmemory.cnt_wr[4] +
             redmule_tb.i_dummy_dmemory.cnt_wr[5] +
             redmule_tb.i_dummy_dmemory.cnt_wr[6] +
             redmule_tb.i_dummy_dmemory.cnt_wr[7] +
             redmule_tb.i_dummy_dmemory.cnt_wr[8];

    $display("[TB] - cnt_rd=%-8d", cnt_rd);
    $display("[TB] - cnt_wr=%-8d", cnt_wr);
    if (perf_enable) begin
      real busy_ratio;
      busy_ratio = (perf_total_cycles != 0) ?
                   (100.0 * real'(perf_busy_cycles) / real'(perf_total_cycles)) : 0.0;
      $display("[PERF] total cycles    : %0d", perf_total_cycles);
      $display("[PERF] busy cycles     : %0d", perf_busy_cycles);
      $display("[PERF] busy ratio      : %0.2f %%", busy_ratio);
      $display("[PERF] MX blocks dec   : %0d", perf_decoder_blocks);
      $display("[PERF] MX blocks enc   : %0d", perf_encoder_blocks);
      $display("[PERF] X stream done   : %0d", x_stream_done_count);
      $display("[PERF] W stream done   : %0d", w_stream_done_count);
      $display("[PERF] Z stream done   : %0d", z_stream_done_count);
    end
    if(errors != 0) begin
      $display("[TB] - Fail!");
      $error("[TB] - errors=%08x", errors);
    end else begin
      $display("[TB] - Success!");
      $display("[TB] - errors=%08x", errors);
    end
    $finish;
  end

  // MX Encoder Output Capture for Verification
  integer mx_fp16_file, mx_fp8_file, mx_exp_file;
  initial begin
    mx_fp16_file = $fopen("mx_encoder_fp16_inputs.txt", "w");
    mx_fp8_file  = $fopen("mx_encoder_fp8_outputs.txt", "w");
    mx_exp_file  = $fopen("mx_encoder_exponents.txt", "w");
  end

  // Capture FP16 inputs when FIFO reads
  always @(posedge clk_i) begin
    if (i_dut.i_redmule_top.fifo_valid && i_dut.i_redmule_top.fifo_pop) begin
      $fwrite(mx_fp16_file, "%h\n", i_dut.i_redmule_top.fifo_data_out);
    end
  end

  // Capture FP8 outputs when encoder produces valid data
  always @(posedge clk_i) begin
    if (i_dut.i_redmule_top.mx_val_valid && i_dut.i_redmule_top.mx_val_ready) begin
      $fwrite(mx_fp8_file, "%h\n", i_dut.i_redmule_top.mx_val_data);
    end
  end

  // Capture shared exponents
  always @(posedge clk_i) begin
    if (i_dut.i_redmule_top.mx_exp_valid && i_dut.i_redmule_top.mx_exp_ready) begin
      $fwrite(mx_exp_file, "%h\n", i_dut.i_redmule_top.mx_exp_data);
    end
  end

  final begin
    $fclose(mx_fp16_file);
    $fclose(mx_fp8_file);
    $fclose(mx_exp_file);
        // Add after simulation ends (near the end of the testbench)
    $display("[TB DEBUG] Memory at y_inp (0x1c0103dc):");
    for (int i = 0; i < 8; i++) begin
      $display("  [%0d]: 0x%08x", i, i_dummy_dmemory.memory[(32'h1c0103dc - 32'h1c010000)/4 + i]);
    end

    $display("[TB DEBUG] Memory at z_oup (check address):");
    // Adjust address based on where z_oup actually is
    $display("[TB] - MX encoder outputs written to mx_encoder_*.txt");
  end

  // always_ff @(posedge clk_i or negedge rst_ni) begin
  //   if (!rst_ni) begin
  //     mx_x_exp_idx <= 0;
  //     mx_w_exp_idx <= 0;
  //   end else begin
  //     // Increment X index only on successful handshake
  //     if (mx_enable && x_mx_exp_stream.valid && x_mx_exp_stream.ready) begin
  //       mx_x_exp_idx <= mx_x_exp_idx + 1;
  //       //$display("[TB][X_EXP] Handshake: idx=%0d data=0x%08x", mx_x_exp_idx, mx_x_exp_mem[mx_x_exp_idx]);
  //     end

  //     // Increment W index only on successful handshake
  //     if (mx_enable && w_mx_exp_stream.valid && w_mx_exp_stream.ready) begin
  //       mx_w_exp_idx <= mx_w_exp_idx + 1;
  //       //$display("[TB][W_EXP] Handshake: idx=%0d data=0x%08x", mx_w_exp_idx, mx_w_exp_mem[mx_w_exp_idx]);
  //     end
  //   end
  // end

endmodule // redmule_tb
